module ForwardingUnit (
  input [3:0] src1, src2, wb_dest, mem_dest,
  input wb_wb_en, mem_wb_en,
  output [1:0] sel_src1, sel_src2
  );

  assign sel_src1 = (mem_wb_en && mem_dest == src1) ? 2'b01 :
                    (wb_wb_en && wb_dest == src1) ? 2'b10 : 2'b00;


  assign sel_src2 = (mem_wb_en && mem_dest == src2) ? 2'b01 :
                    (wb_wb_en && wb_dest == src2) ? 2'b10 : 2'b00;



endmodule